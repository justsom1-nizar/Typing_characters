----------------------------------------------------------------------------------
-- 8x16 Font ROM
-- Converts ASCII character codes to pixel patterns
-- Each character is 8 pixels wide, 16 pixels tall
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.typing_characters_pkg.all;
 
entity font_rom is
    port(
        clk         : in std_logic;
        char_code   : in std_logic_vector(7 downto 0);  -- ASCII code (0-255)
        row         : in integer range 0 to LETTER_HEIGHT;          -- Which row of character (0-15)
        pixel_row   : out std_logic_vector(7 downto 0)  -- 8 pixels for this row
    );
end font_rom;

architecture Behavioral of font_rom is
    
    -- Font data type: array[character][row] = 8 pixels
    type font_row_t is array(0 to 15) of std_logic_vector(7 downto 0);
    type font_rom_t is array(0 to 255) of font_row_t;
    
    -- Font data: IBM VGA style 8x16 font
    -- Each row: MSB (bit 7) is leftmost pixel, LSB (bit 0) is rightmost
    -- '1' = pixel on (foreground), '0' = pixel off (background)
    constant FONT_DATA : font_rom_t := (
        
        -- 0x00-0x1F: Control characters (show as blank or special symbols)
        0 to 31 => (others => x"00"),
        
        -- 0x20: Space
        16#20# => (
            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x21: !
        16#21# => (
            x"00", x"00", x"18", x"18", x"18", x"18", x"18", x"18",
            x"18", x"18", x"00", x"18", x"18", x"00", x"00", x"00"
        ),
        
        -- 0x22: "
        16#22# => (
            x"00", x"66", x"66", x"66", x"24", x"00", x"00", x"00",
            x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x30: 0
        16#30# => (
            x"00", x"00", x"3C", x"66", x"66", x"6E", x"76", x"66",
            x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x31: 1
        16#31# => (
            x"00", x"00", x"18", x"38", x"18", x"18", x"18", x"18",
            x"18", x"18", x"7E", x"00", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x32: 2
        16#32# => (
            x"00", x"00", x"3C", x"66", x"66", x"06", x"0C", x"18",
            x"30", x"60", x"7E", x"00", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x33: 3
        16#33# => (
            x"00", x"00", x"3C", x"66", x"06", x"06", x"1C", x"06",
            x"06", x"66", x"3C", x"00", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x34: 4
        16#34# => (
            x"00", x"00", x"0C", x"1C", x"2C", x"4C", x"4C", x"7E",
            x"0C", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x35: 5
        16#35# => (
            x"00", x"00", x"7E", x"60", x"60", x"7C", x"06", x"06",
            x"06", x"66", x"3C", x"00", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x36: 6
        16#36# => (
            x"00", x"00", x"1C", x"30", x"60", x"7C", x"66", x"66",
            x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x37: 7
        16#37# => (
            x"00", x"00", x"7E", x"06", x"06", x"0C", x"0C", x"18",
            x"18", x"18", x"18", x"00", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x38: 8
        16#38# => (
            x"00", x"00", x"3C", x"66", x"66", x"66", x"3C", x"66",
            x"66", x"66", x"3C", x"00", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x39: 9
        16#39# => (
            x"00", x"00", x"3C", x"66", x"66", x"66", x"3E", x"06",
            x"06", x"0C", x"38", x"00", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x41: A
        16#41# => (
            x"00", x"00", x"18", x"18", x"24", x"24", x"42", x"42",
            x"7E", x"42", x"42", x"42", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x42: B
        16#42# => (
            x"00", x"00", x"7C", x"42", x"42", x"42", x"7C", x"42",
            x"42", x"42", x"42", x"7C", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x43: C
        16#43# => (
            x"00", x"00", x"3C", x"42", x"42", x"40", x"40", x"40",
            x"40", x"42", x"42", x"3C", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x44: D
        16#44# => (
            x"00", x"00", x"78", x"44", x"42", x"42", x"42", x"42",
            x"42", x"42", x"44", x"78", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x45: E
        16#45# => (
            x"00", x"00", x"7E", x"40", x"40", x"40", x"7C", x"40",
            x"40", x"40", x"40", x"7E", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x46: F
        16#46# => (
            x"00", x"00", x"7E", x"40", x"40", x"40", x"7C", x"40",
            x"40", x"40", x"40", x"40", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x47: G
        16#47# => (
            x"00", x"00", x"3C", x"42", x"42", x"40", x"40", x"4E",
            x"42", x"42", x"46", x"3A", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x48: H
        16#48# => (
            x"00", x"00", x"42", x"42", x"42", x"42", x"7E", x"42",
            x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x49: I
        16#49# => (
            x"00", x"00", x"3C", x"18", x"18", x"18", x"18", x"18",
            x"18", x"18", x"18", x"3C", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x4A: J
        16#4A# => (
            x"00", x"00", x"1E", x"0C", x"0C", x"0C", x"0C", x"0C",
            x"0C", x"4C", x"4C", x"38", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x4B: K
        16#4B# => (
            x"00", x"00", x"42", x"44", x"48", x"50", x"60", x"50",
            x"48", x"44", x"42", x"42", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x4C: L
        16#4C# => (
            x"00", x"00", x"40", x"40", x"40", x"40", x"40", x"40",
            x"40", x"40", x"40", x"7E", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x4D: M
        16#4D# => (
            x"00", x"00", x"42", x"42", x"66", x"66", x"5A", x"5A",
            x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x4E: N
        16#4E# => (
            x"00", x"00", x"42", x"42", x"62", x"52", x"4A", x"46",
            x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x4F: O
        16#4F# => (
            x"00", x"00", x"3C", x"42", x"42", x"42", x"42", x"42",
            x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x50: P
        16#50# => (
            x"00", x"00", x"7C", x"42", x"42", x"42", x"7C", x"40",
            x"40", x"40", x"40", x"40", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x51: Q
        16#51# => (
            x"00", x"00", x"3C", x"42", x"42", x"42", x"42", x"42",
            x"42", x"4A", x"44", x"3A", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x52: R
        16#52# => (
            x"00", x"00", x"7C", x"42", x"42", x"42", x"7C", x"50",
            x"48", x"44", x"42", x"42", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x53: S
        16#53# => (
            x"00", x"00", x"3C", x"42", x"40", x"40", x"3C", x"02",
            x"02", x"02", x"42", x"3C", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x54: T
        16#54# => (
            x"00", x"00", x"7E", x"18", x"18", x"18", x"18", x"18",
            x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x55: U
        16#55# => (
            x"00", x"00", x"42", x"42", x"42", x"42", x"42", x"42",
            x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x56: V
        16#56# => (
            x"00", x"00", x"42", x"42", x"42", x"42", x"42", x"42",
            x"42", x"24", x"24", x"18", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x57: W
        16#57# => (
            x"00", x"00", x"42", x"42", x"42", x"42", x"5A", x"5A",
            x"5A", x"66", x"66", x"42", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x58: X
        16#58# => (
            x"00", x"00", x"42", x"42", x"24", x"24", x"18", x"18",
            x"24", x"24", x"42", x"42", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x59: Y
        16#59# => (
            x"00", x"00", x"42", x"42", x"42", x"24", x"24", x"18",
            x"18", x"18", x"18", x"18", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x5A: Z
        16#5A# => (
            x"00", x"00", x"7E", x"02", x"04", x"08", x"10", x"10",
            x"20", x"40", x"40", x"7E", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x61: a (lowercase)
        16#61# => (
            x"00", x"00", x"00", x"00", x"00", x"3C", x"02", x"3E",
            x"42", x"42", x"46", x"3A", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x62: b (lowercase)
        16#62# => (
            x"00", x"00", x"40", x"40", x"40", x"5C", x"62", x"42",
            x"42", x"42", x"62", x"5C", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x63: c (lowercase)
        16#63# => (
            x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"40",
            x"40", x"40", x"42", x"3C", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x64: d (lowercase)
        16#64# => (
            x"00", x"00", x"02", x"02", x"02", x"3A", x"46", x"42",
            x"42", x"42", x"46", x"3A", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x65: e (lowercase)
        16#65# => (
            x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"42",
            x"7E", x"40", x"40", x"3C", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x66: f (lowercase)
        16#66# => (
            x"00", x"00", x"0E", x"10", x"10", x"10", x"7C", x"10",
            x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x67: g (lowercase)
        16#67# => (
            x"00", x"00", x"00", x"00", x"00", x"3A", x"46", x"42",
            x"42", x"46", x"3A", x"02", x"42", x"3C", x"00", x"00"
        ),
        
        -- 0x68: h (lowercase)
        16#68# => (
            x"00", x"00", x"40", x"40", x"40", x"5C", x"62", x"42",
            x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x69: i (lowercase)
        16#69# => (
            x"00", x"00", x"18", x"18", x"00", x"38", x"18", x"18",
            x"18", x"18", x"18", x"3C", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x6A: j (lowercase)
        16#6A# => (
            x"00", x"00", x"0C", x"0C", x"00", x"1C", x"0C", x"0C",
            x"0C", x"0C", x"0C", x"0C", x"4C", x"38", x"00", x"00"
        ),
        
        -- 0x6B: k (lowercase)
        16#6B# => (
            x"00", x"00", x"40", x"40", x"40", x"44", x"48", x"50",
            x"60", x"50", x"48", x"44", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x6C: l (lowercase)
        16#6C# => (
            x"00", x"00", x"38", x"18", x"18", x"18", x"18", x"18",
            x"18", x"18", x"18", x"3C", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x6D: m (lowercase)
        16#6D# => (
            x"00", x"00", x"00", x"00", x"00", x"76", x"49", x"49",
            x"49", x"49", x"49", x"49", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x6E: n (lowercase)
        16#6E# => (
            x"00", x"00", x"00", x"00", x"00", x"5C", x"62", x"42",
            x"42", x"42", x"42", x"42", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x6F: o (lowercase)
        16#6F# => (
            x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"42",
            x"42", x"42", x"42", x"3C", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x70: p (lowercase)
        16#70# => (
            x"00", x"00", x"00", x"00", x"00", x"5C", x"62", x"42",
            x"42", x"62", x"5C", x"40", x"40", x"40", x"00", x"00"
        ),
        
        -- 0x71: q (lowercase)
        16#71# => (
            x"00", x"00", x"00", x"00", x"00", x"3A", x"46", x"42",
            x"42", x"46", x"3A", x"02", x"02", x"02", x"00", x"00"
        ),
        
        -- 0x72: r (lowercase)
        16#72# => (
            x"00", x"00", x"00", x"00", x"00", x"5C", x"62", x"40",
            x"40", x"40", x"40", x"40", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x73: s (lowercase)
        16#73# => (
            x"00", x"00", x"00", x"00", x"00", x"3C", x"42", x"40",
            x"3C", x"02", x"42", x"3C", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x74: t (lowercase)
        16#74# => (
            x"00", x"00", x"00", x"10", x"10", x"7C", x"10", x"10",
            x"10", x"10", x"10", x"0E", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x75: u (lowercase)
        16#75# => (
            x"00", x"00", x"00", x"00", x"00", x"42", x"42", x"42",
            x"42", x"42", x"46", x"3A", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x76: v (lowercase)
        16#76# => (
            x"00", x"00", x"00", x"00", x"00", x"42", x"42", x"42",
            x"42", x"24", x"24", x"18", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x77: w (lowercase)
        16#77# => (
            x"00", x"00", x"00", x"00", x"00", x"42", x"42", x"5A",
            x"5A", x"5A", x"66", x"42", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x78: x (lowercase)
        16#78# => (
            x"00", x"00", x"00", x"00", x"00", x"42", x"24", x"18",
            x"18", x"18", x"24", x"42", x"00", x"00", x"00", x"00"
        ),
        
        -- 0x79: y (lowercase)
        16#79# => (
            x"00", x"00", x"00", x"00", x"00", x"42", x"42", x"42",
            x"42", x"46", x"3A", x"02", x"42", x"3C", x"00", x"00"
        ),
        
        -- 0x7A: z (lowercase)
        16#7A# => (
            x"00", x"00", x"00", x"00", x"00", x"7E", x"04", x"08",
            x"10", x"20", x"40", x"7E", x"00", x"00", x"00", x"00"
        ),
        
        -- Fill remaining characters with blank
        others => (others => x"00")
    );
    
begin
    
    -- Synchronous read
    process(clk)
    begin
        if rising_edge(clk) then
            pixel_row <= FONT_DATA(to_integer(unsigned(char_code)))(row);
        end if;
    end process;
    
end Behavioral;